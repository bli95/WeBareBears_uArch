library verilog;
use verilog.vl_types.all;
entity dcache_ctrlr_sv_unit is
end dcache_ctrlr_sv_unit;
