library verilog;
use verilog.vl_types.all;
entity dcache_phys_mainpc_tb is
end dcache_phys_mainpc_tb;
