library verilog;
use verilog.vl_types.all;
entity VCarray_sv_unit is
end VCarray_sv_unit;
