library verilog;
use verilog.vl_types.all;
entity victim_cache_sv_unit is
end victim_cache_sv_unit;
