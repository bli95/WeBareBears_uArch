library verilog;
use verilog.vl_types.all;
entity mainpc_tb is
end mainpc_tb;
