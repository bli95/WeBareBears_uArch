library verilog;
use verilog.vl_types.all;
entity arbiter is
end arbiter;
