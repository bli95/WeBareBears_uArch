library verilog;
use verilog.vl_types.all;
entity adj_add_pc_sv_unit is
end adj_add_pc_sv_unit;
