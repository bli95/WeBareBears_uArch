library verilog;
use verilog.vl_types.all;
entity LRUarray_sv_unit is
end LRUarray_sv_unit;
