library verilog;
use verilog.vl_types.all;
entity pcmux_ctrlr_sv_unit is
end pcmux_ctrlr_sv_unit;
