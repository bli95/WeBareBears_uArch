library verilog;
use verilog.vl_types.all;
entity VC_LRU_stack_sv_unit is
end VC_LRU_stack_sv_unit;
