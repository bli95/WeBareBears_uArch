library verilog;
use verilog.vl_types.all;
entity mainpc is
end mainpc;
