library verilog;
use verilog.vl_types.all;
entity extend_128_sv_unit is
end extend_128_sv_unit;
