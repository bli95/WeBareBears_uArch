library verilog;
use verilog.vl_types.all;
entity performance_counters_sv_unit is
end performance_counters_sv_unit;
