library verilog;
use verilog.vl_types.all;
entity cpu_rwmod_sv_unit is
end cpu_rwmod_sv_unit;
