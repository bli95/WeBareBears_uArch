library verilog;
use verilog.vl_types.all;
entity cache is
    port(
        level           : in     vl_logic
    );
end cache;
