library verilog;
use verilog.vl_types.all;
entity VC_datapath_sv_unit is
end VC_datapath_sv_unit;
