library verilog;
use verilog.vl_types.all;
entity lc3mask_sv_unit is
end lc3mask_sv_unit;
