library verilog;
use verilog.vl_types.all;
entity write_buffer_sv_unit is
end write_buffer_sv_unit;
