library verilog;
use verilog.vl_types.all;
entity pipeline_sv_unit is
end pipeline_sv_unit;
