library verilog;
use verilog.vl_types.all;
entity BR_array_sv_unit is
end BR_array_sv_unit;
