library verilog;
use verilog.vl_types.all;
entity extract_16_sv_unit is
end extract_16_sv_unit;
