library verilog;
use verilog.vl_types.all;
entity ext_sv_unit is
end ext_sv_unit;
