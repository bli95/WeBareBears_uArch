library verilog;
use verilog.vl_types.all;
entity VC_control_sv_unit is
end VC_control_sv_unit;
