library verilog;
use verilog.vl_types.all;
entity VC_LRUarray_sv_unit is
end VC_LRUarray_sv_unit;
