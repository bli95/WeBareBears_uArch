library verilog;
use verilog.vl_types.all;
entity full_mainpc_tb is
end full_mainpc_tb;
