library verilog;
use verilog.vl_types.all;
entity L2array_sv_unit is
end L2array_sv_unit;
