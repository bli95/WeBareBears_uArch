library verilog;
use verilog.vl_types.all;
entity magic_memory_dual_port is
end magic_memory_dual_port;
