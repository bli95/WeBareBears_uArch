library verilog;
use verilog.vl_types.all;
entity LRU_stack_sv_unit is
end LRU_stack_sv_unit;
