library verilog;
use verilog.vl_types.all;
entity fwd_unit_sv_unit is
end fwd_unit_sv_unit;
