library verilog;
use verilog.vl_types.all;
entity cccomp_sv_unit is
end cccomp_sv_unit;
