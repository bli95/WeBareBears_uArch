library verilog;
use verilog.vl_types.all;
entity sel_bytes_sv_unit is
end sel_bytes_sv_unit;
